/**********************************************************************************************************************
 *  FILE DESCRIPTION
 *  -------------------------------------------------------------------------------------------------------------------
 *  File:         sync_fifo_defines.sv
 *
 *  Description:  
 * 
 *********************************************************************************************************************/

  `ifndef SYNC_FIFO_DEFINES
    `define SYNC_FIFO_DEFINES

    `ifndef FIFO_WIDTH
      `define FIFO_WIDTH    8
    `endif

    `ifndef FIFO_DEPTH
      `define FIFO_DEPTH    8
    `endif 

    `ifndef FIFO_PTR_WIDTH
      `define FIFO_PTR_WIDTH $clog2(`FIFO_DEPTH)
    `endif 
  `endif

/**********************************************************************************************************************
*  END OF FILE: sync_fifo_defines.sv
*********************************************************************************************************************/